package pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"


	`include "seq_item.sv"
	`include "sequence.sv"
	`include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "environment.sv"
	`include "test.sv"

endpackage:pkg
